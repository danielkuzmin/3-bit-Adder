`include full_adder.v

module adder_3bits

(
	input [2:0] a, b,
	input cin,
	output [2:0] sum,
	output co
);



endmodule
